// Copyright 2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Author: Tim Fischer <fischeti@iis.ee.ethz.ch>

`include "axi/assign.svh"
`include "axi/typedef.svh"
`include "tcdm_interface/typedef.svh"

module cluster_tile
  import floo_pkg::*;
  import floo_picobello_noc_pkg::*;
  import snitch_cluster_pkg::*;
  import picobello_pkg::*;
(
  input  logic                                    clk_i,
  input  logic                                    rst_ni,
  input  logic                                    test_enable_i,
  input  logic                                    tile_clk_en_i,
  input  logic                                    tile_rst_ni,
  input  logic                                    clk_rst_bypass_i,
  // Cluster ports
  input  logic                      [NrCores-1:0] debug_req_i,
  input  logic                      [NrCores-1:0] meip_i,
  input  logic                      [NrCores-1:0] mtip_i,
  input  logic                      [NrCores-1:0] msip_i,
  input  logic                      [        9:0] hart_base_id_i,
  input  snitch_cluster_pkg::addr_t               cluster_base_addr_i,
  input  snitch_cluster_pkg::addr_t               cluster_base_offset_i,
  // Chimney ports
  input  id_t                                     id_i,
  // Router ports
  output floo_req_t                 [ West:North] floo_req_o,
  input  floo_rsp_t                 [ West:North] floo_rsp_i,
  output floo_wide_t                [ West:North] floo_wide_o,
  input  floo_req_t                 [ West:North] floo_req_i,
  output floo_rsp_t                 [ West:North] floo_rsp_o,
  input  floo_wide_t                [ West:North] floo_wide_i
);

  /// TODO(lleone): Offload typedef to be generated by Floogen or removed form
  /// the hardware after more optimization
  typedef logic[AxiCfgW.DataWidth-1:0] RdDataWide_t;
  typedef logic[AxiCfgN.DataWidth-1:0] RdDataNarrow_t;


  // Tile-specific reset and clock signals
  logic                                 tile_clk;
  logic                                 tile_rst_n;

  ////////////////////
  // Snitch Cluster //
  ////////////////////

  snitch_cluster_pkg::narrow_in_req_t   cluster_narrow_in_req;
  snitch_cluster_pkg::narrow_in_resp_t  cluster_narrow_in_rsp;
  snitch_cluster_pkg::narrow_out_req_t  cluster_narrow_out_req;
  snitch_cluster_pkg::narrow_out_resp_t cluster_narrow_out_rsp;
  snitch_cluster_pkg::wide_out_req_t    cluster_wide_out_req;
  snitch_cluster_pkg::wide_out_resp_t   cluster_wide_out_rsp;
  snitch_cluster_pkg::wide_in_req_t     cluster_wide_in_req;
  snitch_cluster_pkg::wide_in_resp_t    cluster_wide_in_rsp;

  snitch_cluster_pkg::narrow_out_req_t  cluster_narrow_ext_req;
  snitch_cluster_pkg::narrow_out_resp_t cluster_narrow_ext_rsp;
  snitch_cluster_pkg::tcdm_dma_req_t    cluster_tcdm_ext_req_aligned;
  snitch_cluster_pkg::tcdm_dma_req_t    cluster_tcdm_ext_req_misaligned;
  snitch_cluster_pkg::tcdm_dma_rsp_t    cluster_tcdm_ext_rsp_aligned;
  snitch_cluster_pkg::tcdm_dma_rsp_t    cluster_tcdm_ext_rsp_misaligned;

  localparam int unsigned HWPECtrlAddrWidth = 32;
  localparam int unsigned HWPECtrlDataWidth = 32;
  typedef logic [HWPECtrlAddrWidth-1:0] addr_hwpe_ctrl_t;
  typedef logic [HWPECtrlDataWidth-1:0] data_hwpe_ctrl_t;
  typedef logic [3:0] strb_hwpe_ctrl_t;

  `AXI_TYPEDEF_ALL(cluster_narrow_out_dw_conv, snitch_cluster_pkg::addr_t,
                   snitch_cluster_pkg::narrow_out_id_t, data_hwpe_ctrl_t, strb_hwpe_ctrl_t,
                   snitch_cluster_pkg::user_narrow_t)

  cluster_narrow_out_dw_conv_req_t cluster_narrow_out_dw_conv_req, cluster_narrow_out_cut_req;
  cluster_narrow_out_dw_conv_resp_t cluster_narrow_out_dw_conv_rsp, cluster_narrow_out_cut_rsp;

  `TCDM_TYPEDEF_ALL(hwpectrl, addr_hwpe_ctrl_t, data_hwpe_ctrl_t, strb_hwpe_ctrl_t, logic)

  hwpectrl_req_t               hwpectrl_req;
  hwpectrl_rsp_t               hwpectrl_rsp;

  logic          [NrCores-1:0] mxip;


  ////////////////////////
  // Wide FPU Reduction //
  ////////////////////////

  // Snitch cluster DCA interface
  snitch_cluster_pkg::dca_req_t offload_dca_req, offload_dca_req_cut;
  snitch_cluster_pkg::dca_rsp_t offload_dca_rsp, offload_dca_rsp_cut;

  // Signals to connect the NW router to the wide parser
  RdDataWide_t [1:0]  offload_wide_req_operand;
  collect_op_e        offload_wide_req_operation;
  logic               offload_wide_req_valid;
  logic               offload_wide_req_ready;
  RdDataWide_t        offload_wide_resp_data;
  logic               offload_wide_resp_valid;
  logic               offload_wide_resp_ready;

  // Parse the Wide request from the reouter to the one from the snitch cluster!
  // TODO(raroth): possible to remove this decode from the picobello repo and move it inside the
  //       FlooNoC repo. Currently the Decode used for the ALU is directly inside the floo_alu.sv
  //       file. Maybe do the same for the FPU
  if(EnWideOffloadReduction) begin : gen_wide_offload_reduction
    // Connect the DCA Request
    assign offload_dca_req.q_valid = offload_wide_req_valid;
    assign offload_wide_req_ready = offload_dca_rsp.q_ready;

    // Parse the FPU Request
    always_comb begin
      // Init default values
      offload_dca_req.q.operands = '0;

      // Set default Values
      offload_dca_req.q.src_fmt = fpnew_pkg::FP64;
      offload_dca_req.q.dst_fmt = fpnew_pkg::FP64;
      offload_dca_req.q.int_fmt = fpnew_pkg::INT64;
      offload_dca_req.q.vectorial_op = 1'b0;
      offload_dca_req.q.op_mod = 1'b0;
      offload_dca_req.q.rnd_mode = fpnew_pkg::RNE;
      offload_dca_req.q.op = fpnew_pkg::ADD;

      // Define the operation we want to execute on the FPU
      unique casez (offload_wide_req_operation)
        (floo_pkg::F_Add) : begin
          offload_dca_req.q.op = fpnew_pkg::ADD;
          offload_dca_req.q.operands[0] = '0;
          offload_dca_req.q.operands[1] = offload_wide_req_operand[0];
          offload_dca_req.q.operands[2] = offload_wide_req_operand[1];
        end
        (floo_pkg::F_Mul) : begin
          offload_dca_req.q.op = fpnew_pkg::MUL;
          offload_dca_req.q.operands[0] = offload_wide_req_operand[0];
          offload_dca_req.q.operands[1] = offload_wide_req_operand[1];
          offload_dca_req.q.operands[2] = '0;
        end
        (floo_pkg::F_Max) : begin
          offload_dca_req.q.op = fpnew_pkg::MINMAX;
          offload_dca_req.q.rnd_mode = fpnew_pkg::RNE;
          offload_dca_req.q.operands[0] = offload_wide_req_operand[0];
          offload_dca_req.q.operands[1] = offload_wide_req_operand[1];
          offload_dca_req.q.operands[2] = '0;
        end
        (floo_pkg::F_Min) : begin
          offload_dca_req.q.op = fpnew_pkg::MINMAX;
          offload_dca_req.q.rnd_mode = fpnew_pkg::RTZ;
          offload_dca_req.q.operands[0] = offload_wide_req_operand[0];
          offload_dca_req.q.operands[1] = offload_wide_req_operand[1];
          offload_dca_req.q.operands[2] = '0;
        end
        default : begin
          offload_dca_req.q.op = fpnew_pkg::ADD;
          offload_dca_req.q.operands[0] = '0;
          offload_dca_req.q.operands[1] = '0;
          offload_dca_req.q.operands[2] = '0;
        end
      endcase
    end

    // TODO(raroth): move these spill register inside FlooNoC and make them configurable.
    // Insert a reqrsp-cut to avoid timing violations
    generic_reqrsp_cut #(
      .req_chan_t (snitch_cluster_pkg::dca_req_chan_t),
      .rsp_chan_t (snitch_cluster_pkg::dca_rsp_chan_t),
      .BypassReq  (1'b0),
      .BypassRsp  (1'b0)
    ) i_dca_router_cut (
      .clk_i          (clk_i),
      .rst_ni         (rst_ni),
      .slv_req_i      (offload_dca_req),
      .slv_rsp_o      (offload_dca_rsp),
      .mst_req_o      (offload_dca_req_cut),
      .mst_rsp_i      (offload_dca_rsp_cut)
    );
    // Connect the Response
    assign offload_wide_resp_valid = offload_dca_rsp.p_valid;
    assign offload_dca_req.p_ready = offload_wide_resp_ready;
    assign offload_wide_resp_data = offload_dca_rsp.p.result;

  // No Wide Reduction supported
  end else begin : gen_no_wide_reduction
    assign offload_dca_req_cut = '0;
    assign offload_dca_rsp = '0;
    assign offload_wide_req_ready = '0;
    assign offload_wide_resp_data = '0;
    assign offload_wide_resp_valid = '0;
  end

  // TODO(lleone): Add teh narrow ALU reduction unit and connections here


  snitch_cluster_wrapper i_cluster (
    .clk_i            (tile_clk),
    .rst_ni           (tile_rst_n),
    .debug_req_i,
    .meip_i,
    .mtip_i,
    .msip_i,
    .hart_base_id_i,
    .cluster_base_addr_i,
    .cluster_base_offset_i,
    .mxip_i           (mxip),
    .clk_d2_bypass_i  ('0),
    .sram_cfgs_i      ('0),
    .narrow_in_req_i  (cluster_narrow_in_req),
    .narrow_in_resp_o (cluster_narrow_in_rsp),
    .narrow_out_req_o (cluster_narrow_out_req),
    .narrow_out_resp_i(cluster_narrow_out_rsp),
    .wide_out_req_o   (cluster_wide_out_req),
    .wide_out_resp_i  (cluster_wide_out_rsp),
    .wide_in_req_i    (cluster_wide_in_req),
    .wide_in_resp_o   (cluster_wide_in_rsp),
    .narrow_ext_req_o (cluster_narrow_ext_req),
    .narrow_ext_resp_i(cluster_narrow_ext_rsp),
    .tcdm_ext_req_i   (cluster_tcdm_ext_req_aligned),
    .tcdm_ext_resp_o  (cluster_tcdm_ext_rsp_aligned),
    .dca_req_i        (offload_dca_req_cut),
    .dca_rsp_o        (offload_dca_rsp_cut)
  );

  // Convert narrow AXI's 64 bit DW down to 32
  axi_dw_converter #(
    .AxiMaxReads        (1),
    .AxiSlvPortDataWidth(snitch_cluster_pkg::NarrowDataWidth),
    .AxiMstPortDataWidth(HWPECtrlDataWidth),
    .AxiAddrWidth       (snitch_cluster_pkg::AddrWidth),
    .AxiIdWidth         (snitch_cluster_pkg::NarrowIdWidthOut),
    .aw_chan_t          (snitch_cluster_pkg::narrow_out_aw_chan_t),
    .mst_w_chan_t       (cluster_narrow_out_dw_conv_w_chan_t),
    .slv_w_chan_t       (snitch_cluster_pkg::narrow_out_w_chan_t),
    .b_chan_t           (snitch_cluster_pkg::narrow_out_b_chan_t),
    .ar_chan_t          (snitch_cluster_pkg::narrow_out_ar_chan_t),
    .mst_r_chan_t       (cluster_narrow_out_dw_conv_r_chan_t),
    .slv_r_chan_t       (snitch_cluster_pkg::narrow_out_r_chan_t),
    .axi_mst_req_t      (cluster_narrow_out_dw_conv_req_t),
    .axi_mst_resp_t     (cluster_narrow_out_dw_conv_resp_t),
    .axi_slv_req_t      (snitch_cluster_pkg::narrow_out_req_t),
    .axi_slv_resp_t     (snitch_cluster_pkg::narrow_out_resp_t)
  ) i_axi_dw_hwpe (
    .clk_i     (tile_clk),
    .rst_ni    (tile_rst_n),
    .slv_req_i (cluster_narrow_ext_req),
    .slv_resp_o(cluster_narrow_ext_rsp),
    .mst_req_o (cluster_narrow_out_dw_conv_req),
    .mst_resp_i(cluster_narrow_out_dw_conv_rsp)
  );

  axi_cut #(
    .Bypass    (0),
    .aw_chan_t (snitch_cluster_pkg::narrow_out_aw_chan_t),
    .w_chan_t  (cluster_narrow_out_dw_conv_w_chan_t),
    .b_chan_t  (snitch_cluster_pkg::narrow_out_b_chan_t),
    .ar_chan_t (snitch_cluster_pkg::narrow_out_ar_chan_t),
    .r_chan_t  (cluster_narrow_out_dw_conv_r_chan_t),
    .axi_req_t (cluster_narrow_out_dw_conv_req_t),
    .axi_resp_t(cluster_narrow_out_dw_conv_resp_t)
  ) i_cut_ext_narrow_slv (
    .clk_i     (tile_clk),
    .rst_ni    (tile_rst_n),
    .slv_req_i (cluster_narrow_out_dw_conv_req),
    .slv_resp_o(cluster_narrow_out_dw_conv_rsp),
    .mst_req_o (cluster_narrow_out_cut_req),
    .mst_resp_i(cluster_narrow_out_cut_rsp)
  );

  axi_to_tcdm #(
    .axi_req_t (cluster_narrow_out_dw_conv_req_t),
    .axi_rsp_t (cluster_narrow_out_dw_conv_resp_t),
    .tcdm_req_t(hwpectrl_req_t),
    .tcdm_rsp_t(hwpectrl_rsp_t),
    .IdWidth   (snitch_cluster_pkg::NarrowIdWidthOut),
    .AddrWidth (HWPECtrlAddrWidth),
    .DataWidth (HWPECtrlDataWidth)
  ) i_axi_to_hwpe_ctrl (
    .clk_i     (tile_clk),
    .rst_ni    (tile_rst_n),
    .axi_req_i (cluster_narrow_out_cut_req),
    .axi_rsp_o (cluster_narrow_out_cut_rsp),
    .tcdm_req_o(hwpectrl_req),
    .tcdm_rsp_i(hwpectrl_rsp)
  );

  snitch_tcdm_aligner #(
    .tcdm_req_t   (snitch_cluster_pkg::tcdm_dma_req_t),
    .tcdm_rsp_t   (snitch_cluster_pkg::tcdm_dma_rsp_t),
    .DataWidth    (snitch_cluster_pkg::WideDataWidth),
    .TCDMDataWidth(snitch_cluster_pkg::NarrowDataWidth),
    .AddrWidth    (snitch_cluster_pkg::TcdmAddrWidth)
  ) i_snitch_tcdm_aligner (
    .clk_i                (tile_clk),
    .rst_ni               (tile_rst_n),
    .tcdm_req_misaligned_i(cluster_tcdm_ext_req_misaligned),
    .tcdm_req_aligned_o   (cluster_tcdm_ext_req_aligned),
    .tcdm_rsp_aligned_i   (cluster_tcdm_ext_rsp_aligned),
    .tcdm_rsp_misaligned_o(cluster_tcdm_ext_rsp_misaligned)
  );

  snitch_hwpe_subsystem #(
    .tcdm_req_t   (snitch_cluster_pkg::tcdm_dma_req_t),
    .tcdm_rsp_t   (snitch_cluster_pkg::tcdm_dma_rsp_t),
    .periph_req_t (hwpectrl_req_t),
    .periph_rsp_t (hwpectrl_rsp_t),
    .HwpeDataWidth(snitch_cluster_pkg::WideDataWidth),
    .IdWidth      (snitch_cluster_pkg::NarrowIdWidthOut),
    .NrCores      (NrCores),
    .TCDMDataWidth(snitch_cluster_pkg::NarrowDataWidth)
  ) i_snitch_hwpe_subsystem (
    .clk_i          (tile_clk),
    .rst_ni         (tile_rst_n),
    .test_mode_i    (1'b0),
    .tcdm_req_o     (cluster_tcdm_ext_req_misaligned),
    .tcdm_rsp_i     (cluster_tcdm_ext_rsp_misaligned),
    .hwpe_ctrl_req_i(hwpectrl_req),
    .hwpe_ctrl_rsp_o(hwpectrl_rsp),
    .hwpe_evt_o     (mxip)
  );

  ////////////
  // Router //
  ////////////

  typedef struct packed {
    logic [1:0] valid;
    logic [1:0] ready;
    floo_wide_chan_t [1:0] wide;
  } floo_wide_double_t;

  floo_req_t [Eject:North] router_floo_req_out, router_floo_req_in;
  floo_rsp_t [Eject:North] router_floo_rsp_out, router_floo_rsp_in;
  floo_wide_double_t [Eject:North] router_floo_wide_out;
  floo_wide_t [Eject:North] router_floo_wide_in;

  floo_nw_router_v2 #(
    .AxiCfgN     (AxiCfgN),
    .AxiCfgW     (AxiCfgW),
    .RouteAlgo   (RouteCfg.RouteAlgo),
    .EnMultiCast (RouteCfg.EnMultiCast),
    .EnParallelReduction      (EnParallelReduction),
    .EnOffloadWideReduction   (EnWideOffloadReduction),
    .EnOffloadNarrowReduction (EnNarrowOffloadReduction),
    .EnDecoupledRW (1'b1),
    .NoLoopback  (1'b0),
    .NumRoutes   (5),
    .InFifoDepth (2),
    .OutFifoDepth(2),
    .id_t        (id_t),
    .hdr_t       (hdr_t),
    .floo_req_t  (floo_req_t),
    .floo_rsp_t  (floo_rsp_t),
    .floo_wide_t (floo_wide_t),
    .floo_wide_out_t (floo_wide_double_t),
    .RdWideOperation_t        (floo_pkg::collect_op_e),
    .RdNarrowOperation_t      (floo_pkg::collect_op_e),
    .RdWideData_t             (RdDataWide_t),
    .RdNarrowData_t           (RdDataNarrow_t),
    .RdWideCfg                (WideReductionCfg),
    .RdNarrowCfg              (NarrowReductionCfg),
    .RdRespCfg                (ResponseReductionCfg)
  ) i_router (
    .clk_i,
    .rst_ni,
    .test_enable_i,
    .id_i,
    .id_route_map_i('0),
    .floo_req_i    (router_floo_req_in),
    .floo_rsp_o    (router_floo_rsp_out),
    .floo_req_o    (router_floo_req_out),
    .floo_rsp_i    (router_floo_rsp_in),
    .floo_wide_i   (router_floo_wide_in),
    .floo_wide_o   (router_floo_wide_out),
    // Wide Reduction offload port
    .offload_wide_req_op_o          (offload_wide_req_operation),
    .offload_wide_req_operand1_o    (offload_wide_req_operand[0]),
    .offload_wide_req_operand2_o    (offload_wide_req_operand[1]),
    .offload_wide_req_valid_o       (offload_wide_req_valid),
    .offload_wide_req_ready_i       (offload_wide_req_ready),
    .offload_wide_resp_result_i     (offload_wide_resp_data),
    .offload_wide_resp_valid_i      (offload_wide_resp_valid),
    .offload_wide_resp_ready_o      (offload_wide_resp_ready),
    // Narrow Reduction offload port
    .offload_narrow_req_op_o        (),
    .offload_narrow_req_operand1_o  (),
    .offload_narrow_req_operand2_o  (),
    .offload_narrow_req_valid_o     (),
    .offload_narrow_req_ready_i     ('0),
    .offload_narrow_resp_result_i   ('0),
    .offload_narrow_resp_valid_i    ('0),
    .offload_narrow_resp_ready_o    ()
  );

  assign floo_req_o                      = router_floo_req_out[West:North];
  assign router_floo_req_in[West:North]  = floo_req_i;
  assign floo_rsp_o                      = router_floo_rsp_out[West:North];
  assign router_floo_rsp_in[West:North]  = floo_rsp_i;
  // Only the local port uses both physical channels. Other outputs use only the lower.
  for (genvar i = North; i <= West; i++) begin : gen_floo_wide_o
    assign floo_wide_o[i].valid = router_floo_wide_out[i].valid;
    assign floo_wide_o[i].ready = router_floo_wide_out[i].ready;
    assign floo_wide_o[i].wide = router_floo_wide_out[i].wide[0];
  end
  assign router_floo_wide_in[West:North] = floo_wide_i;

  /////////////
  // Chimney //
  /////////////

  floo_nw_chimney_v2 #(
    .AxiCfgN             (floo_picobello_noc_pkg::AxiCfgN),
    .AxiCfgW             (floo_picobello_noc_pkg::AxiCfgW),
    .ChimneyCfgN         (floo_pkg::ChimneyDefaultCfg),
    .ChimneyCfgW         (floo_pkg::ChimneyDefaultCfg),
    .RouteCfg            (floo_picobello_noc_pkg::RouteCfg),
    .AtopSupport         (1'b1),
    .EnDecoupledRW       (1'b1),
    .MaxAtomicTxns       (1),
    .Sam                 (picobello_pkg::SamMcast),
    .id_t                (floo_picobello_noc_pkg::id_t),
    .rob_idx_t           (floo_picobello_noc_pkg::rob_idx_t),
    .hdr_t               (floo_picobello_noc_pkg::hdr_t),
    .sam_rule_t          (picobello_pkg::sam_multicast_rule_t),
    .sam_idx_t           (picobello_pkg::sam_idx_t),
    .mask_sel_t          (picobello_pkg::mask_sel_t),
    .axi_narrow_in_req_t (snitch_cluster_pkg::narrow_out_req_t),
    .axi_narrow_in_rsp_t (snitch_cluster_pkg::narrow_out_resp_t),
    .axi_narrow_out_req_t(snitch_cluster_pkg::narrow_in_req_t),
    .axi_narrow_out_rsp_t(snitch_cluster_pkg::narrow_in_resp_t),
    .axi_wide_in_req_t   (snitch_cluster_pkg::wide_out_req_t),
    .axi_wide_in_rsp_t   (snitch_cluster_pkg::wide_out_resp_t),
    .axi_wide_out_req_t  (snitch_cluster_pkg::wide_in_req_t),
    .axi_wide_out_rsp_t  (snitch_cluster_pkg::wide_in_resp_t),
    .floo_req_t          (floo_picobello_noc_pkg::floo_req_t),
    .floo_rsp_t          (floo_picobello_noc_pkg::floo_rsp_t),
    .floo_wide_t         (floo_picobello_noc_pkg::floo_wide_t),
    .floo_wide_in_t         (floo_wide_double_t),
    .sram_cfg_t          (snitch_cluster_pkg::sram_cfg_t),
    .user_narrow_struct_t         (picobello_pkg::collective_narrow_user_t),
    .user_wide_struct_t           (picobello_pkg::collective_wide_user_t)
  ) i_chimney (
    .clk_i               (tile_clk),
    .rst_ni              (tile_rst_n),
    .test_enable_i,
    .id_i,
    .route_table_i       ('0),
    .sram_cfg_i          ('0),
    .axi_narrow_in_req_i (cluster_narrow_out_req),
    .axi_narrow_in_rsp_o (cluster_narrow_out_rsp),
    .axi_narrow_out_req_o(cluster_narrow_in_req),
    .axi_narrow_out_rsp_i(cluster_narrow_in_rsp),
    .axi_wide_in_req_i   (cluster_wide_out_req),
    .axi_wide_in_rsp_o   (cluster_wide_out_rsp),
    .axi_wide_out_req_o  (cluster_wide_in_req),
    .axi_wide_out_rsp_i  (cluster_wide_in_rsp),
    .floo_req_o          (router_floo_req_in[Eject]),
    .floo_rsp_o          (router_floo_rsp_in[Eject]),
    .floo_wide_o         (router_floo_wide_in[Eject]),
    .floo_req_i          (router_floo_req_out[Eject]),
    .floo_rsp_i          (router_floo_rsp_out[Eject]),
    .floo_wide_i         (router_floo_wide_out[Eject])
  );

  //////////////////////////
  // Clock Gating & Reset //
  //////////////////////////

  tc_clk_gating i_tc_clk_gating_cluster (
    .clk_i,
    .en_i     (tile_clk_en_i),
    .test_en_i(clk_rst_bypass_i),
    .clk_o    (tile_clk)
  );

`ifdef TARGET_XILINX
  // Using clk cells makes Vivado flag the reset as a clock tree
  assign tile_rst_n = (clk_rst_bypass_i) ? rst_ni : tile_rst_ni;
`else
  tc_clk_mux2 i_tc_reset_mux (
    .clk0_i   (tile_rst_ni),
    .clk1_i   (rst_ni),
    .clk_sel_i(clk_rst_bypass_i),
    .clk_o    (tile_rst_n)
  );
`endif



endmodule
