// Copyright 2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Author: Tim Fischer <fischeti@iis.ee.ethz.ch>

`include "axi/assign.svh"

module sparta_tile
  import floo_pkg::*;
  import floo_picobello_noc_pkg::*;
  import picobello_pkg::*;
(
  input  logic clk_i,
  input  logic rst_ni,
  input  logic test_enable_i,
  // Cluster ports
  input  logic [snitch_cluster_pkg::NrCores-1:0] debug_req_i,
  input  logic [snitch_cluster_pkg::NrCores-1:0] meip_i,
  input  logic [snitch_cluster_pkg::NrCores-1:0] mtip_i,
  input  logic [snitch_cluster_pkg::NrCores-1:0] msip_i,
  input  logic [9:0]                             hart_base_id_i,
  input  snitch_cluster_pkg::addr_t              cluster_base_addr_i,
  // Chimney ports
  input  id_t id_i,
  // Router ports
  output floo_req_t [West:North]    floo_req_o,
  input  floo_rsp_t [West:North]    floo_rsp_i,
  output floo_wide_t [West:North]   floo_wide_o,
  input  floo_req_t [West:North]    floo_req_i,
  output floo_rsp_t [West:North]    floo_rsp_o,
  input  floo_wide_t [West:North]   floo_wide_i
);

  snitch_cluster_pkg::narrow_in_req_t   cluster_narrow_in_req;
  snitch_cluster_pkg::narrow_in_resp_t  cluster_narrow_in_rsp;
  snitch_cluster_pkg::narrow_out_req_t  cluster_narrow_out_req;
  snitch_cluster_pkg::narrow_out_resp_t cluster_narrow_out_rsp;
  snitch_cluster_pkg::wide_out_req_t    cluster_wide_out_req;
  snitch_cluster_pkg::wide_out_resp_t   cluster_wide_out_rsp;
  snitch_cluster_pkg::wide_in_req_t     cluster_wide_in_req;
  snitch_cluster_pkg::wide_in_resp_t    cluster_wide_in_rsp;

  snitch_cluster_wrapper i_cluster (
    .clk_i                ( clk_i                   ),
    .rst_ni               ( rst_ni                  ),
    .debug_req_i          ( debug_req_i             ),
    .meip_i               ( meip_i                  ),
    .mtip_i               ( mtip_i                  ),
    .msip_i               ( msip_i                  ),
    .hart_base_id_i       ( hart_base_id_i          ),
    .cluster_base_addr_i  ( cluster_base_addr_i     ),
    .clk_d2_bypass_i      ( '0                      ),
    .sram_cfgs_i          ( '0                      ),
    .narrow_in_req_i      ( cluster_narrow_in_req   ),
    .narrow_in_resp_o     ( cluster_narrow_in_rsp   ),
    .narrow_out_req_o     ( cluster_narrow_out_req  ),
    .narrow_out_resp_i    ( cluster_narrow_out_rsp  ),
    .wide_out_req_o       ( cluster_wide_out_req    ),
    .wide_out_resp_i      ( cluster_wide_out_rsp    ),
    .wide_in_req_i        ( cluster_wide_in_req     ),
    .wide_in_resp_o       ( cluster_wide_in_rsp     )
  );

  floo_picobello_noc_pkg::axi_narrow_in_req_t  chimney_narrow_in_req;
  floo_picobello_noc_pkg::axi_narrow_in_rsp_t  chimney_narrow_in_rsp;
  floo_picobello_noc_pkg::axi_narrow_out_req_t chimney_narrow_out_req;
  floo_picobello_noc_pkg::axi_narrow_out_rsp_t chimney_narrow_out_rsp;
  floo_picobello_noc_pkg::axi_wide_out_req_t   chimney_wide_out_req;
  floo_picobello_noc_pkg::axi_wide_out_rsp_t   chimney_wide_out_rsp;
  floo_picobello_noc_pkg::axi_wide_in_req_t    chimney_wide_in_req;
  floo_picobello_noc_pkg::axi_wide_in_rsp_t    chimney_wide_in_rsp;

  `AXI_ASSIGN_REQ_STRUCT(cluster_narrow_in_req, chimney_narrow_out_req);
  `AXI_ASSIGN_RESP_STRUCT(chimney_narrow_out_rsp, cluster_narrow_in_rsp);
  `AXI_ASSIGN_REQ_STRUCT(chimney_narrow_in_req, cluster_narrow_out_req);
  `AXI_ASSIGN_RESP_STRUCT(cluster_narrow_out_rsp, chimney_narrow_in_rsp);
  `AXI_ASSIGN_REQ_STRUCT(cluster_wide_in_req, chimney_wide_out_req);
  `AXI_ASSIGN_RESP_STRUCT(chimney_wide_out_rsp, cluster_wide_in_rsp);
  `AXI_ASSIGN_REQ_STRUCT(chimney_wide_in_req, cluster_wide_out_req);
  `AXI_ASSIGN_RESP_STRUCT(cluster_wide_out_rsp, chimney_wide_in_rsp);

  floo_req_t  [Eject:North] router_floo_req_out, router_floo_req_in;
  floo_rsp_t  [Eject:North] router_floo_rsp_out, router_floo_rsp_in;
  floo_wide_t [Eject:North] router_floo_wide_out, router_floo_wide_in;

  floo_nw_chimney #(
    .AxiCfgN              ( floo_picobello_noc_pkg::AxiCfgN              ),
    .AxiCfgW              ( floo_picobello_noc_pkg::AxiCfgW              ),
    .ChimneyCfgN          ( floo_pkg::ChimneyDefaultCfg                  ),
    .ChimneyCfgW          ( floo_pkg::ChimneyDefaultCfg                  ),
    .RouteCfg             ( floo_picobello_noc_pkg::RouteCfg             ),
    .AtopSupport          ( 1'b1                                         ),
    .MaxAtomicTxns        ( 1                                            ),
    .Sam                  ( floo_picobello_noc_pkg::Sam                  ),
    .id_t                 ( floo_picobello_noc_pkg::id_t                 ),
    .rob_idx_t            ( floo_picobello_noc_pkg::rob_idx_t            ),
    .hdr_t                ( floo_picobello_noc_pkg::hdr_t                ),
    .sam_rule_t           ( floo_picobello_noc_pkg::sam_rule_t           ),
    .axi_narrow_in_req_t  ( floo_picobello_noc_pkg::axi_narrow_in_req_t  ),
    .axi_narrow_in_rsp_t  ( floo_picobello_noc_pkg::axi_narrow_in_rsp_t  ),
    .axi_narrow_out_req_t ( floo_picobello_noc_pkg::axi_narrow_out_req_t ),
    .axi_narrow_out_rsp_t ( floo_picobello_noc_pkg::axi_narrow_out_rsp_t ),
    .axi_wide_in_req_t    ( floo_picobello_noc_pkg::axi_wide_in_req_t    ),
    .axi_wide_in_rsp_t    ( floo_picobello_noc_pkg::axi_wide_in_rsp_t    ),
    .axi_wide_out_req_t   ( floo_picobello_noc_pkg::axi_wide_out_req_t   ),
    .axi_wide_out_rsp_t   ( floo_picobello_noc_pkg::axi_wide_out_rsp_t   ),
    .floo_req_t           ( floo_picobello_noc_pkg::floo_req_t           ),
    .floo_rsp_t           ( floo_picobello_noc_pkg::floo_rsp_t           ),
    .floo_wide_t          ( floo_picobello_noc_pkg::floo_wide_t          ),
    .sram_cfg_t           ( snitch_cluster_pkg::sram_cfg_t               )
  ) i_chimney (
    .clk_i,
    .rst_ni,
    .test_enable_i,
    .id_i,
    .route_table_i        ( '0                          ),
    .sram_cfg_i           ( '0                          ),
    .axi_narrow_in_req_i  ( chimney_narrow_in_req       ),
    .axi_narrow_in_rsp_o  ( chimney_narrow_in_rsp       ),
    .axi_narrow_out_req_o ( chimney_narrow_out_req      ),
    .axi_narrow_out_rsp_i ( chimney_narrow_out_rsp      ),
    .axi_wide_in_req_i    ( chimney_wide_in_req         ),
    .axi_wide_in_rsp_o    ( chimney_wide_in_rsp         ),
    .axi_wide_out_req_o   ( chimney_wide_out_req        ),
    .axi_wide_out_rsp_i   ( chimney_wide_out_rsp        ),
    .floo_req_o           ( router_floo_req_in[Eject]   ),
    .floo_rsp_o           ( router_floo_rsp_in[Eject]   ),
    .floo_wide_o          ( router_floo_wide_in[Eject]  ),
    .floo_req_i           ( router_floo_req_out[Eject]  ),
    .floo_rsp_i           ( router_floo_rsp_out[Eject]  ),
    .floo_wide_i          ( router_floo_wide_out[Eject] )
  );

  floo_nw_router #(
    .AxiCfgN      ( AxiCfgN             ),
    .AxiCfgW      ( AxiCfgW             ),
    .RouteAlgo    ( RouteCfg.RouteAlgo  ),
    .NumRoutes    ( 5                   ),
    .InFifoDepth  ( 2                   ),
    .OutFifoDepth ( 2                   ),
    .id_t         ( id_t                ),
    .hdr_t        ( hdr_t               ),
    .floo_req_t   ( floo_req_t          ),
    .floo_rsp_t   ( floo_rsp_t          ),
    .floo_wide_t  ( floo_wide_t         )
  ) i_router (
    .clk_i,
    .rst_ni,
    .test_enable_i,
    .id_i,
    .id_route_map_i ( '0                    ),
    .floo_req_i     ( router_floo_req_in    ),
    .floo_rsp_o     ( router_floo_rsp_out   ),
    .floo_req_o     ( router_floo_req_out   ),
    .floo_rsp_i     ( router_floo_rsp_in    ),
    .floo_wide_i    ( router_floo_wide_in   ),
    .floo_wide_o    ( router_floo_wide_out  )
  );

  assign floo_req_o = router_floo_req_out[West:North];
  assign router_floo_req_in[West:North] = floo_req_i;
  assign floo_rsp_o = router_floo_rsp_out[West:North];
  assign router_floo_rsp_in[West:North] = floo_rsp_i;
  assign floo_wide_o = router_floo_wide_out[West:North];
  assign router_floo_wide_in[West:North] = floo_wide_i;

endmodule
